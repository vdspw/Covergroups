/*this is an FSM for which we are ging to write an example to demonstrate usage of illegal bins */

module state_mach(
input rst,clk,
input din,
output logic dout
);
 
parameter s0 = 2'b00;
parameter s1 = 2'b01;
parameter s2 = 2'b10;
  
  reg [1:0] state, next_state;  ///00-11 is the actual range but we dont want the design to reach 11 (3) , if it does its operation is wrong (ERROR).
 
/////////////Reset Logic
always_ff@(posedge clk)
begin
if(rst == 1'b1)
state <= s0;
else
state <= next_state;
end
 
///////////////Next state Decoder Logic
always_comb
begin
  case(state)
s0: begin
if(din == 1'b1)
next_state = s1;
else
next_state = s0;
end
 
s1: begin
if(din == 1'b1)
next_state = s2;
else
next_state = s1;
end
  
s2: begin
if(din == 1'b1)
next_state = s0;
else
next_state = s2;
end  
 
default : next_state = s0;
endcase
end
 
///////////////Output Logic
 
always_comb
begin
case(state)
s0: dout = 1'b0;
s1: dout = 1'b0;
s2: dout = 1'b1;  
default : dout = 1'b0;
endcase
end
 
 
 
endmodule
/////////////////////////////////////////////////////////////////////////////////////////////////


//////////////////////// TB code
/* to flag the state 3(11) as an ERROR we must include it in the illegal_bins
this is done in both state and next_state */


module tb;
  
  reg clk = 0;
  reg reset = 0;
  reg din = 0;
  wire dout;
  
 
 state_mach dut (reset,clk,din, dout);
  
 always #5 clk = ~clk;
  
  initial begin
    reset = 1;
    #30;
    reset = 0;
    #40;
    din = 1;
  end
 
 
  covergroup c;
    option.per_instance = 1;
    
    coverpoint dut.state iff (!reset){
    
      bins fsmstate[] = {0,1,2}; //states for which covergae will be calculated.
      illegal_bins unused_state = {3};
    }
    
    coverpoint dut.next_state iff (!reset){
    
      bins fsmstate[] = {0,1,2};//states for which covergae will be calculated.
      illegal_bins unused_state = {3};
    }
    
  endgroup
  
    c ci;
    
    initial begin
      ci = new();
      forever begin
        @(posedge clk);
        ci.sample();
      end
    end
 
  
  
  
  
 initial begin
    $dumpfile("dump.vcd"); 
    $dumpvars;
    #300;
    $finish();
  end
  
 
endmodule
