/* Ignore bins part 2 */ 
/* value A can range from 0 to 255 ,we are condiering values 1 to 100 only ,
we want to ignore tha value 23,45,67,89,93 */

module tb;
  
  reg [7:0] a;
  integer i = 0;
 
  
  covergroup c;
    option.per_instance = 1;
    
    coverpoint a {
      bins value_a[] = {[1:100]};
      ignore_bins unused_a = {23,45,67,89,93};    
    }
    
    
    
  endgroup
  
  
  
  
  
 
  
 
  c ci;
 
  initial begin
     ci = new();
    
    
    
    for (i = 0; i <40; i++) begin
      a = $urandom();
      ci.sample();
      #10;
    end
    
    
  end
  
  
  
  
  initial begin
    $dumpfile("dump.vcd"); 
    $dumpvars;
    #400;
    $finish();
  end
  
 
 
 
 
endmodule
